// FPGA Design Control FSM Module
// Henry Heathwood
// hheathwood@hmc.edu
// 11/18/24

module control_FSM(input logic [7:0] value, logic [4:0] paramOut, logic SPIDone, logic dataDone, logic clk, logic reset,
					output logic dataReady, logic RSin, logic RWin, logic [7:0] dataIn);
					
					
endmodule